module array_divider_6bit(
    input [5:0] A, B,
    );

    


endmodule